../../lib/reconos_defs.vhd