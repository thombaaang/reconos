../hls/mbox/solution1/syn/vhdl/top.vhd