../hls/mbox/solution1/syn/vhdl/FIFO_top_queue_get_V_V.vhd