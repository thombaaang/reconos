../../../../reconos_defs.vhd