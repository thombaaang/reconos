../../lib/thread/reconos_thread_vhdl.vhd