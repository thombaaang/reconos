../../lib/thread/reconos_calls_vhdl.vhd