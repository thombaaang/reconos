../hls/mbox/solution1/syn/vhdl/FIFO_top_queue_put_V_V.vhd