../sim_thread_14.7/reconos_testbench.vhd