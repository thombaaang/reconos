../hls/mbox/solution1/syn/vhdl/FIFO_top_mbox_V_V.vhd